import ovm_pkg::*;
import bdb_tb_transactions_pkg::*;

module  bdb_tb_comparator (
  ref tlm_fifo #(bdb_result) actual_result_fifo,
  ref tlm_fifo #(bdb_result) predicted_result_fifo
);
	
	bdb_result actual_result;
  bdb_result predicted_result;
  string m;
  string message;
		
	task run;
	  
	  $sformat(m, "%m");
	  
	  forever begin
	   
	    actual_result_fifo.get(actual_result);
	    predicted_result_fifo.get(predicted_result);
	   
	     $sformat(message, "Predicted: %s   Actual: %s",
	       predicted_result.convert2string, actual_result.convert2string);
	   
      if (actual_result.comp(predicted_result))
        ovm_top.ovm_report_info(m, message, 300);
      else 
        ovm_top.ovm_report_error(m, message, 200);
	   
	   end  
	 
	endtask
	 
endmodule

