`define FIFO_WIDTH 4
