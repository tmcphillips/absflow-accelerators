
module reverse_complement_demo (
	input			wire					clock_100m
);

	
 complement_soc u0 (
	  .clk_clk 			(clock_100m)
 );

endmodule

